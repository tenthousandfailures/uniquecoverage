package TB0_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "TB0_env.sv"
`include "TB0_test.sv"

endpackage // TB0_pkg
    
